module fpgaTop(
input clk
);
endmodule 
module RAM_1PORT ();

integer i;
always begin
end
endmodule